`include "pcie_defs.vh"
`include "nif_common_defs.vh"

////////////////////////////////////////
//{{{ SLAVE INTERFACE
////////////////////////////////////////
`define NIF_SLAVE_ADDRESS_WIDTH									64
`define NIF_SLAVE_CS_WIDTH										4
`define NIF_SLAVE_BE_WIDTH										16
`define NIF_SLAVE_DATA_WIDTH									128

`define NIF_SLAVE_IF_CMD_WIDTH									128

`define NIF_SLAVE_IF_CMD_TYPE_WIDTH								4
`define NIF_SLAVE_IF_CMD_TYPE_LOW								0
`define NIF_SLAVE_IF_CMD_TYPE_HIGH								(`NIF_SLAVE_IF_CMD_TYPE_LOW + `NIF_SLAVE_IF_CMD_TYPE_WIDTH - 1)
`define NIF_SLAVE_IF_CMD_TYPE_FIELD								(`NIF_SLAVE_IF_CMD_TYPE_HIGH):(`NIF_SLAVE_IF_CMD_TYPE_LOW)

`define NIF_SLAVE_IF_CMD_BURST_SIZE_WIDTH						16
`define NIF_SLAVE_IF_CMD_BURST_SIZE_LOW							(`NIF_SLAVE_IF_CMD_TYPE_HIGH + 1)
`define NIF_SLAVE_IF_CMD_BURST_SIZE_HIGH						(`NIF_SLAVE_IF_CMD_BURST_SIZE_LOW + `NIF_SLAVE_IF_CMD_BURST_SIZE_WIDTH - 1)
`define NIF_SLAVE_IF_CMD_BURST_SIZE_FIELD						(`NIF_SLAVE_IF_CMD_BURST_SIZE_HIGH):(`NIF_SLAVE_IF_CMD_BURST_SIZE_LOW)

`define NIF_SLAVE_IF_CMD_BURST_STRIDE_WIDTH						16
`define NIF_SLAVE_IF_CMD_BURST_STRIDE_LOW						(`NIF_SLAVE_IF_CMD_BURST_SIZE_HIGH + 1)
`define NIF_SLAVE_IF_CMD_BURST_STRIDE_HIGH						(`NIF_SLAVE_IF_CMD_BURST_STRIDE_LOW + `NIF_SLAVE_IF_CMD_BURST_STRIDE_WIDTH - 1)
`define NIF_SLAVE_IF_CMD_BURST_STRIDE_FIELD						(`NIF_SLAVE_IF_CMD_BURST_STRIDE_HIGH):(`NIF_SLAVE_IF_CMD_BURST_STRIDE_LOW)

`define NIF_SLAVE_IF_CMD_LENGTH_WIDTH							20
`define NIF_SLAVE_IF_CMD_LENGTH_LOW								(`NIF_SLAVE_IF_CMD_BURST_STRIDE_HIGH + 1)
`define NIF_SLAVE_IF_CMD_LENGTH_HIGH							(`NIF_SLAVE_IF_CMD_LENGTH_LOW + `NIF_SLAVE_IF_CMD_LENGTH_WIDTH - 1)
`define NIF_SLAVE_IF_CMD_LENGTH_FIELD							(`NIF_SLAVE_IF_CMD_LENGTH_HIGH):(`NIF_SLAVE_IF_CMD_LENGTH_LOW)

`define NIF_SLAVE_IF_CMD_TRANSACTION_OPTIONS_WIDTH				4
`define NIF_SLAVE_IF_CMD_TRANSACTION_OPTIONS_LOW				(`NIF_SLAVE_IF_CMD_LENGTH_HIGH + 1)
`define	NIF_SLAVE_IF_CMD_TRANSACTION_OPTIONS_HIGH				(`NIF_SLAVE_IF_CMD_TRANSACTION_OPTIONS_LOW + `NIF_SLAVE_IF_CMD_TRANSACTION_OPTIONS_WIDTH - 1)
`define NIF_SLAVE_IF_CMD_TRANSACTION_OPTIONS_FIELD				(`NIF_SLAVE_IF_CMD_TRANSACTION_OPTIONS_HIGH):(`NIF_SLAVE_IF_CMD_TRANSACTION_OPTIONS_LOW)

`define NIF_SLAVE_IF_CMD_SLAVE_SELECT_FLAG						(`NIF_SLAVE_IF_CMD_TRANSACTION_OPTIONS_HIGH + 1)
`define NIF_SLAVE_IF_CMD_EOF_FLAG								(`NIF_SLAVE_IF_CMD_SLAVE_SELECT_FLAG + 1)

`define NIF_SLAVE_IF_CMD_CS_WIDTH								2
`define NIF_SLAVE_IF_CMD_CS_LOW									(`NIF_SLAVE_IF_CMD_EOF_FLAG + 1)
`define NIF_SLAVE_IF_CMD_CS_HIGH								(`NIF_SLAVE_IF_CMD_CS_LOW + `NIF_SLAVE_IF_CMD_CS_WIDTH - 1)
`define NIF_SLAVE_IF_CMD_CS_FIELD								(`NIF_SLAVE_IF_CMD_CS_HIGH):(`NIF_SLAVE_IF_CMD_CS_LOW)

`define NIF_SLAVE_IF_CMD_ADDRESS_WIDTH							64
`define NIF_SLAVE_IF_CMD_ADDRESS_LOW							64
`define NIF_SLAVE_IF_CMD_ADDRESS_HIGH							(`NIF_SLAVE_IF_CMD_ADDRESS_LOW + `NIF_SLAVE_IF_CMD_ADDRESS_WIDTH - 1)
`define NIF_SLAVE_IF_CMD_ADDRESS_FIELD							(`NIF_SLAVE_IF_CMD_ADDRESS_HIGH):(`NIF_SLAVE_IF_CMD_ADDRESS_LOW)

`define NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_ADDRESS_WIDTH		(`NIF_SLAVE_IF_CMD_ADDRESS_WIDTH)
`define NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_ADDRESS_LOW		0
`define NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_ADDRESS_HIGH		(`NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_ADDRESS_LOW + `NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_ADDRESS_WIDTH - 1)
`define NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_ADDRESS_FIELD		(`NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_ADDRESS_HIGH):(`NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_ADDRESS_LOW)

`define NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_CHIPSELECT_WIDTH	(`NIF_SLAVE_CS_WIDTH)
`define NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_CHIPSELECT_LOW		(`NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_ADDRESS_HIGH + 1)
`define NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_CHIPSELECT_HIGH	(`NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_ADDRESS_HIGH + `NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_CHIPSELECT_WIDTH - 1)
`define NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_CHIPSELECT_FIELD	(`NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_CHIPSELECT_HIGH):(`NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_CHIPSELECT_LOW)

`define NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_WIDTH				(`NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_ADDRESS_WIDTH + `NIF_SLAVE_IF_ADDRESS_LOOKUP_RESPONSE_CHIPSELECT_WIDTH)

// Definition of Slave Interface Command Types
`define NIF_SLAVE_IF_CMD_TYPE_1D_READ	4'd0
`define NIF_SLAVE_IF_CMD_TYPE_1D_WRITE	4'd1

// Definition of Maximum Read Length from Slave Interface
`define DMA_SLAVE_READ_MAX_BYTE					2048
`define LOG2_DMA_SLAVE_READ_MAX_BYTE			11

////////////////////////////////////////
//}}} SLAVE INTERFACE
////////////////////////////////////////



////////////////////////////////////////
//{{{ Static System Memory Space Allocation
////////////////////////////////////////
// ---------------------------------
// 16 total spaces = 12 system spaces + 4 application spaces
//
// Each system memory has 256 MB memory space.
// Total system memory has 12 x 256 MB + 1024 MB (Reserved Space) = 3072 MB + 1024 MB = 4GB memory space.
// 
//
// Remaining 60 GB out of 64 GB can be dynamically allocated into 4 additional application memory spaces.
// ---------------------------------

`define	NIF_SLAVE_IF_MEM0_BASEADDR		36'h0_0000_0000		// Configuration Handler0
`define NIF_SLAVE_IF_MEM1_BASEADDR		36'h0_1000_0000		// Configuration Handler1
`define NIF_SLAVE_IF_MEM2_BASEADDR		36'h0_2000_0000		// Configuration Handler2
`define NIF_SLAVE_IF_MEM3_BASEADDR		36'h0_3000_0000		// Configuration Handler3
`define NIF_SLAVE_IF_MEM4_BASEADDR		36'h0_4000_0000		// Configuration Handler4
`define NIF_SLAVE_IF_MEM5_BASEADDR		36'h0_5000_0000		// Configuration Handler5
`define NIF_SLAVE_IF_MEM6_BASEADDR		36'h0_6000_0000		// Configuration Handler6
`define NIF_SLAVE_IF_MEM7_BASEADDR		36'h0_7000_0000		// Configuration Handler7
`define NIF_SLAVE_IF_MEM8_BASEADDR		36'h0_8000_0000		// Configuration Packet Egress
`define NIF_SLAVE_IF_MEM9_BASEADDR		36'h0_9000_0000		// Configuration Slave Interface
`define NIF_SLAVE_IF_MEM10_BASEADDR		36'h0_A000_0000		// 
`define NIF_SLAVE_IF_MEM11_BASEADDR		36'h0_B000_0000		//
`define NIF_SLAVE_IF_MEM12_BASEADDR		36'h0_C000_0000		// Application Space0
`define NIF_SLAVE_IF_MEM13_BASEADDR_DEF	36'hF_FFFF_FFFF		// Application Space1 (Default)
`define NIF_SLAVE_IF_MEM14_BASEADDR_DEF	36'hF_FFFF_FFFF		// Application Space2 (Default)
`define NIF_SLAVE_IF_MEM15_BASEADDR_DEF	36'hF_FFFF_FFFF		// Application Space3 (Default)
// Base address of MEM13 ~ MEM15 will be dynamically configured through "Slave Interface Configuration".

////////////////////////////////////////
//}}} Static System Memory Space Allocation
////////////////////////////////////////



////////////////////////////////////////
//{{{ MEMORY REQUEST PACKET FORMAT
////////////////////////////////////////

// ----(Header)-------------------------
// Length		= Always 4DW
// Type, Fmt	= Memory Write 4DW w/data Header
// Tag			= {1'b0, 3'Target Handler ID, 4'Ticket Number}
// ----(Payload)-------------------------
// Req Length, Req Flow
// --------------------------------------

`define	MEMREQ_PAYLOAD_ADDRESS_WIDTH			36
`define	MEMREQ_PAYLOAD_ADDRESS_LOW				0
`define	MEMREQ_PAYLOAD_ADDRESS_HIGH				(`MEMREQ_PAYLOAD_ADDRESS_LOW + `MEMREQ_PAYLOAD_ADDRESS_WIDTH - 1)
`define	MEMREQ_PAYLOAD_ADDRESS_FIELD			(`MEMREQ_PAYLOAD_ADDRESS_HIGH):(`MEMREQ_PAYLOAD_ADDRESS_LOW)

`define MEMREQ_PAYLOAD_LENGTH_WIDTH				36
`define MEMREQ_PAYLOAD_LENGTH_LOW				(`MEMREQ_PAYLOAD_ADDRESS_HIGH + 1)
`define MEMREQ_PAYLOAD_LENGTH_HIGH				(`MEMREQ_PAYLOAD_LENGTH_LOW + `MEMREQ_PAYLOAD_LENGTH_WIDTH - 1)
`define	MEMREQ_PAYLOAD_LENGTH_FIELD				(`MEMREQ_PAYLOAD_LENGTH_HIGH):(`MEMREQ_PAYLOAD_LENGTH_LOW)

`define MEMREQ_PAYLOAD_FLOW_WIDTH				10
`define MEMREQ_PAYLOAD_FLOW_LOW					(`MEMREQ_PAYLOAD_LENGTH_HIGH + 1)
`define MEMREQ_PAYLOAD_FLOW_HIGH				(`MEMREQ_PAYLOAD_FLOW_LOW + `MEMREQ_PAYLOAD_FLOW_WIDTH - 1)
`define	MEMREQ_PAYLOAD_FLOW_FIELD				(`MEMREQ_PAYLOAD_FLOW_HIGH):(`MEMREQ_PAYLOAD_FLOW_LOW)

`define	MEMREQ_PAYLOAD_CONVERGING_FLOW_WIDTH	10
`define	MEMREQ_PAYLOAD_CONVERGING_FLOW_LOW		(`MEMREQ_PAYLOAD_FLOW_HIGH + 1)
`define	MEMREQ_PAYLOAD_CONVERGING_FLOW_HIGH		(`MEMREQ_PAYLOAD_CONVERGING_FLOW_LOW + `MEMREQ_PAYLOAD_CONVERGING_FLOW_WIDTH - 1)
`define	MEMREQ_PAYLOAD_CONVERGING_FLOW_FIELD	(`MEMREQ_PAYLOAD_CONVERGING_FLOW_HIGH):(`MEMREQ_PAYLOAD_CONVERGING_FLOW_LOW)

`define MEMREQ_PAYLOAD_ADDRESS_MSB_WIDTH		28
`define	MEMREQ_PAYLOAD_ADDRESS_MSB_LOW			(`MEMREQ_PAYLOAD_CONVERGING_FLOW_HIGH + 1)
`define	MEMREQ_PAYLOAD_ADDRESS_MSB_HIGH			(`MEMREQ_PAYLOAD_ADDRESS_MSB_LOW + `MEMREQ_PAYLOAD_ADDRESS_MSB_WIDTH - 1)
`define	MEMREQ_PAYLOAD_ADDRESS_MSB_FIELD		(`MEMREQ_PAYLOAD_ADDRESS_MSB_HIGH):(`MEMREQ_PAYLOAD_ADDRESS_MSB_LOW)

`define MEMREQ_PAYLOAD_ADDRESS_EXT_WIDTH	64	


`define MEMREQ_PAYLOAD_RSVD_WIDTH				36

////////////////////////////////////////
//}}} MEMORY REQUEST PACKET FORMAT
////////////////////////////////////////



////////////////////////////////////////
//{{{ EGRESS INTERFACE
////////////////////////////////////////

// ---------------------------------
// Definition of Command Fields
// ---------------------------------
`define	NIF_EGRESS_CMD_COMMAND_WIDTH			6
`define NIF_EGRESS_CMD_COMMAND_LOW				0
`define NIF_EGRESS_CMD_COMMAND_HIGH				(`NIF_EGRESS_CMD_COMMAND_LOW + `NIF_EGRESS_CMD_COMMAND_WIDTH - 1)
`define	NIF_EGRESS_CMD_COMMAND_FIELD			(`NIF_EGRESS_CMD_COMMAND_HIGH):(`NIF_EGRESS_CMD_COMMAND_LOW)

`define	NIF_EGRESS_CMD_FLOW_ID_WIDTH			10
`define NIF_EGRESS_CMD_FLOW_ID_LOW				(`NIF_EGRESS_CMD_COMMAND_HIGH + 1)
`define NIF_EGRESS_CMD_FLOW_ID_HIGH				(`NIF_EGRESS_CMD_FLOW_ID_LOW + `NIF_EGRESS_CMD_FLOW_ID_WIDTH - 1)
`define	NIF_EGRESS_CMD_FLOW_ID_FIELD			(`NIF_EGRESS_CMD_FLOW_ID_HIGH):(`NIF_EGRESS_CMD_FLOW_ID_LOW)

`define	NIF_EGRESS_CMD_DEVICE_ID_WIDTH			16
`define NIF_EGRESS_CMD_DEVICE_ID_LOW 			(`NIF_EGRESS_CMD_FLOW_ID_HIGH + 1)
`define NIF_EGRESS_CMD_DEVICE_ID_HIGH 			(`NIF_EGRESS_CMD_DEVICE_ID_LOW + `NIF_EGRESS_CMD_DEVICE_ID_WIDTH - 1)
`define	NIF_EGRESS_CMD_DEVICE_ID_FIELD			(`NIF_EGRESS_CMD_DEVICE_ID_HIGH):(`NIF_EGRESS_CMD_DEVICE_ID_LOW)

`define	NIF_EGRESS_CMD_ADDRESS_WIDTH			64
`define NIF_EGRESS_CMD_ADDRESS_LOW				(`NIF_EGRESS_CMD_DEVICE_ID_HIGH + 1)
`define NIF_EGRESS_CMD_ADDRESS_HIGH				(`NIF_EGRESS_CMD_ADDRESS_LOW + `NIF_EGRESS_CMD_ADDRESS_WIDTH - 1)
`define	NIF_EGRESS_CMD_ADDRESS_FIELD			(`NIF_EGRESS_CMD_ADDRESS_HIGH):(`NIF_EGRESS_CMD_ADDRESS_LOW)
`define NIF_EGRESS_CMD_ADDRESS_L30_HIGH			(`NIF_EGRESS_CMD_ADDRESS_LOW + 32 - 1 ) 


`define	NIF_EGRESS_CMD_LENGTH_WIDTH				36
`define NIF_EGRESS_CMD_LENGTH_LOW				(`NIF_EGRESS_CMD_ADDRESS_HIGH + 1)
`define NIF_EGRESS_CMD_LENGTH_HIGH				(`NIF_EGRESS_CMD_LENGTH_LOW + `NIF_EGRESS_CMD_LENGTH_WIDTH - 1)
`define	NIF_EGRESS_CMD_LENGTH_FIELD				(`NIF_EGRESS_CMD_LENGTH_HIGH):(`NIF_EGRESS_CMD_LENGTH_LOW)

`define	NIF_EGRESS_CMD_TAG_WIDTH				8
`define NIF_EGRESS_CMD_TAG_LOW					(`NIF_EGRESS_CMD_LENGTH_HIGH + 1)
`define NIF_EGRESS_CMD_TAG_HIGH					(`NIF_EGRESS_CMD_TAG_LOW + `NIF_EGRESS_CMD_TAG_WIDTH - 1)
`define	NIF_EGRESS_CMD_TAG_FIELD				(`NIF_EGRESS_CMD_TAG_HIGH):(`NIF_EGRESS_CMD_TAG_LOW)

`define	NIF_EGRESS_CMD_ERRCODE_WIDTH			7
`define NIF_EGRESS_CMD_ERRCODE_LOW				(`NIF_EGRESS_CMD_TAG_HIGH + 1)
`define NIF_EGRESS_CMD_ERRCODE_HIGH				(`NIF_EGRESS_CMD_ERRCODE_LOW + `NIF_EGRESS_CMD_ERRCODE_WIDTH - 1)
`define	NIF_EGRESS_CMD_ERRCODE_FIELD			(`NIF_EGRESS_CMD_ERRCODE_HIGH):(`NIF_EGRESS_CMD_ERRCODE_LOW)

`define	NIF_EGRESS_CMD_1ST_DW_BE_WIDTH			4
`define NIF_EGRESS_CMD_1ST_DW_BE_LOW			(`NIF_EGRESS_CMD_ERRCODE_HIGH + 1)
`define NIF_EGRESS_CMD_1ST_DW_BE_HIGH			(`NIF_EGRESS_CMD_1ST_DW_BE_LOW + `NIF_EGRESS_CMD_1ST_DW_BE_WIDTH - 1)
`define	NIF_EGRESS_CMD_1ST_DW_BE_FIELD			(`NIF_EGRESS_CMD_1ST_DW_BE_HIGH):(`NIF_EGRESS_CMD_1ST_DW_BE_LOW)

`define	NIF_EGRESS_CMD_LAST_DW_BE_WIDTH			4
`define NIF_EGRESS_CMD_LAST_DW_BE_LOW			(`NIF_EGRESS_CMD_1ST_DW_BE_HIGH + 1)
`define NIF_EGRESS_CMD_LAST_DW_BE_HIGH			(`NIF_EGRESS_CMD_LAST_DW_BE_LOW + `NIF_EGRESS_CMD_LAST_DW_BE_WIDTH - 1)
`define	NIF_EGRESS_CMD_LAST_DW_BE_FIELD			(`NIF_EGRESS_CMD_LAST_DW_BE_HIGH):(`NIF_EGRESS_CMD_LAST_DW_BE_LOW)

`define	NIF_EGRESS_CMD_TRANSACTION_ID_WIDTH		4
`define NIF_EGRESS_CMD_TRANSACTION_ID_LOW		(`NIF_EGRESS_CMD_LAST_DW_BE_HIGH + 1)
`define NIF_EGRESS_CMD_TRANSACTION_ID_HIGH		(`NIF_EGRESS_CMD_TRANSACTION_ID_LOW + `NIF_EGRESS_CMD_TRANSACTION_ID_WIDTH - 1)
`define	NIF_EGRESS_CMD_TRANSACTION_ID_FIELD		(`NIF_EGRESS_CMD_TRANSACTION_ID_HIGH):(`NIF_EGRESS_CMD_TRANSACTION_ID_LOW)

`define	NIF_EGRESS_CMD_RESERVED_FLAG			(`NIF_EGRESS_CMD_TRANSACTION_ID_HIGH + 1)

`define	NIF_EGRESS_CMD_CONVFLOW_ID_WIDTH		10
`define	NIF_EGRESS_CMD_CONVFLOW_ID_LOW			(`NIF_EGRESS_CMD_RESERVED_FLAG + 1)
`define	NIF_EGRESS_CMD_CONVFLOW_ID_HIGH			(`NIF_EGRESS_CMD_CONVFLOW_ID_LOW + `NIF_EGRESS_CMD_CONVFLOW_ID_WIDTH -1)
`define	NIF_EGRESS_CMD_CONVFLOW_ID_FIELD		(`NIF_EGRESS_CMD_CONVFLOW_ID_HIGH):(`NIF_EGRESS_CMD_CONVFLOW_ID_LOW)

// added 9-26-2014

`define NIF_EGRESS_CMD_WIDTH 	(`NIF_EGRESS_CMD_COMMAND_WIDTH	+ 	`NIF_EGRESS_CMD_FLOW_ID_WIDTH + `NIF_EGRESS_CMD_DEVICE_ID_WIDTH + `NIF_EGRESS_CMD_ADDRESS_WIDTH + 	`NIF_EGRESS_CMD_LENGTH_WIDTH + 	`NIF_EGRESS_CMD_TAG_WIDTH + `NIF_EGRESS_CMD_ERRCODE_WIDTH + `NIF_EGRESS_CMD_1ST_DW_BE_WIDTH + `NIF_EGRESS_CMD_LAST_DW_BE_WIDTH + `NIF_EGRESS_CMD_TRANSACTION_ID_WIDTH + `NIF_EGRESS_CMD_CONVFLOW_ID_WIDTH + 1)

`define NIF_EGRESS_ERR_CMD_WIDTH (`NIF_EGRESS_CMD_WIDTH - `NIF_EGRESS_CMD_CONVFLOW_ID_WIDTH)

//Moved to pcie_defs.vh since NIF_SOP is also referencing it..
//`define PCIE_MEM_WRREQ_HEADER_DEFAULT		({32'd0,32'd0,32'd0,1'd0,`PCIE_FMT_FIELD_DEFAULT,`PCIE_TYPE_FIELD_DEFAULT,1'd0,3'd0,4'd0,`PCIE_TD_FIELD_DEFAULT,`PCIE_EP_FIELD_DEFAULT,`PCIE_ATTR_FIELD_DEFAULT,2'd0,10'd0})

// ---------------------------------
// Definition of Command Types
// ---------------------------------
`define NIF_EGRESS_CMD_ERROR						`SYSTEM_FLOW_ID_ERROR
`define NIF_EGRESS_CMD_RSV_REQ_CRITICAL				`SYSTEM_FLOW_ID_RSV_REQ_CRITICAL	
`define NIF_EGRESS_CMD_RSV_REQ_BEST_CHANCE			`SYSTEM_FLOW_ID_RSV_REQ_BEST_CHANCE
`define NIF_EGRESS_CMD_RSV_REQ_BEST_EFFORT			`SYSTEM_FLOW_ID_RSV_REQ_BEST_EFFORT
`define NIF_EGRESS_CMD_WRITE_REQUEST				`SYSTEM_FLOW_ID_WRITE_REQUEST
`define NIF_EGRESS_CMD_WRITE_ACK					`SYSTEM_FLOW_ID_WRITE_ACK
`define	NIF_EGRESS_CMD_WRITE_CANCEL					`SYSTEM_FLOW_ID_WRITE_CANCEL
`define NIF_EGRESS_CMD_WRITE_COMPLETE				`SYSTEM_FLOW_ID_WRITE_COMPLETE
`define NIF_EGRESS_CMD_WRITE_DATA					`SYSTEM_FLOW_ID_WRITE_DATA
`define NIF_EGRESS_CMD_READ_REQUEST					`SYSTEM_FLOW_ID_READ_REQUEST
`define	NIF_EGRESS_CMD_READ_ACK						`SYSTEM_FLOW_ID_READ_ACK
`define	NIF_EGRESS_CMD_READ_START					`SYSTEM_FLOW_ID_READ_START
`define	NIF_EGRESS_CMD_READ_CANCEL					`SYSTEM_FLOW_ID_READ_CANCEL
`define NIF_EGRESS_CMD_READ_COMPLETE				`SYSTEM_FLOW_ID_READ_COMPLETE
`define NIF_EGRESS_CMD_SINGLE_WRITE					`SYSTEM_FLOW_ID_SINGLE_WRITE
`define NIF_EGRESS_CMD_SINGLE_READ					`SYSTEM_FLOW_ID_SINGLE_READ

////////////////////////////////////////
//}}} EGRESS INTERFACE
////////////////////////////////////////


 
////////////////////////////////////////
//{{{ NIF SAP HANDLER STATUS DEFINITION
////////////////////////////////////////

`define NIF_HANDLER_STATUS_IDLE						2'd0
`define NIF_HANDLER_STATUS_BUSY_EXCEPT_ALLOWED		2'd1
`define NIF_HANDLER_STATUS_BUSY_NO_EXCEPTION		2'd2

////////////////////////////////////////
//}}} NIF SAP HANDLER STATUS DEFINITION
////////////////////////////////////////



////////////////////////////////////////
//{{{ NIF SAP ERROR CODE DEFINITION
////////////////////////////////////////

`define	NIF_ERRCODE_NO_ERROR						7'd0
`define NIF_ERRCODE_HANDLER_BUSY					7'd1
`define NIF_ERRCODE_UNEXPECTED_REPLY_FROM_REMOTE	7'd2
`define NIF_ERRCODE_UNSUPPORTED_CMD					7'd3	// Kevin, should we combine this and the bottom one? - Sungho
`define NIF_ERRCODE_UNSUPPORTED_CMD_SLAVE_IF		7'd4
`define NIF_ERRCODE_EGRESS_EARLY_TERMINATION		7'd5
`define NIF_ERRCODE_SLAVE_EARLY_TERMINATION			7'd6
`define NIF_ERRCODE_NO_HANDLER_RESPONSE				7'd7
`define	NIF_ERRCODE_NO_MSG_HANDLER_EXISTS			7'd8
`define	NIF_ERRCODE_NO_ASSOCIATIVE_HANDLER			7'd9
`define NIF_ERRCODE_INVALID_ARGUMENT				7'd10
`define NIF_ERRCODE_TRANSACTION_EARLY_TERMINATION	7'd11
`define NIF_ERRCODE_UNKNOWN_DEVICE_ID				7'd12
////////////////////////////////////////
//}}} NIF SAP ERROR CODE DEFINITION
////////////////////////////////////////



////////////////////////////////////////
//{{{ MASTER INTERFACE
////////////////////////////////////////

// ---------------------------------
// NIF SAP MASTER COMMAND TYPE DEFINITION
// ---------------------------------
`define	NIF_MASTER_CMD_WIDTH						4

`define NIF_MASTER_CMD_WRREQ						4'd0	// Master --> (Remote Device or Local Slave)
`define NIF_MASTER_CMD_RDREQ						4'd1	// (Remote Device or Local Slave) --> Master
`define NIF_MASTER_CMD_WRREQ_DMA					4'd2	// (Local Slave) --> (Remote Slave)
`define NIF_MASTER_CMD_RDREQ_DMA					4'd3	// (Remote Slave) --> (Local Slave)
`define NIF_MASTER_CMD_WRREQ_SINGLE					4'd4	// Master --> (Remote Device or Local Slave) with a small amount of data (less than 4KB)
`define NIF_MASTER_CMD_RDREQ_SINGLE					4'd5	// (Remote Device or Local Slave) --> Master with a small amount of data (less than 4KB)
`define NIF_MASTER_CMD_WRREQ_WINDOW					4'd6	// Master --> (Remote Device or Local Slave) Windowed
`define NIF_MASTER_CMD_RDREQ_WINDOW					4'd7	// (Remote Device or Local Slave) --> Master Windowed
`define NIF_MASTER_CMD_CANCEL						4'd8	// Cancel an active transaction

`define NIF_CMD_VARIANT_NONE						4'd0	// Read/Write no variant
`define NIF_CMD_VARIANT_ALLOCATE_MODIFIED			4'd1	// Read/Write allocate within cache in modified state
`define NIF_CMD_VARIANT_ALLOCATE_SHARED				4'd2	// Read/Write allocate within cache in modified state and transistion to shared state when snooped
`define NIF_CMD_VARIANT_ALLOCATE_RESERVED			4'd3	// Read and create a reservation in the cache
`define NIF_CMD_VARIANT_NO_ALLOCATE					4'd4	// Read/Write no allocate
`define NIF_CMD_VARIANT_NO_ALLOCATE_INJECT			4'd5	// Write no allocate and inject in highest point of coherence

// ---------------------------------
// NIF SAP MASTER COMMAND OPTIONS FIELD DEFINITION
// ---------------------------------
`define NIF_MASTER_CMD_OPTION_LENGTH_WIDTH				36
`define NIF_MASTER_CMD_OPTION_LENGTH_LOW				0
`define NIF_MASTER_CMD_OPTION_LENGTH_HIGH				(`NIF_MASTER_CMD_OPTION_LENGTH_LOW + `NIF_MASTER_CMD_OPTION_LENGTH_WIDTH - 1)
`define	NIF_MASTER_CMD_OPTION_LENGTH_FIELD				(`NIF_MASTER_CMD_OPTION_LENGTH_HIGH):(`NIF_MASTER_CMD_OPTION_LENGTH_LOW)

`define NIF_MASTER_CMD_OPTION_LOCAL_ADDR_WIDTH			36
`define NIF_MASTER_CMD_OPTION_LOCAL_ADDR_LOW			(`NIF_MASTER_CMD_OPTION_LENGTH_HIGH + 1)
`define NIF_MASTER_CMD_OPTION_LOCAL_ADDR_HIGH			(`NIF_MASTER_CMD_OPTION_LOCAL_ADDR_LOW + `NIF_MASTER_CMD_OPTION_LOCAL_ADDR_WIDTH - 1)
`define	NIF_MASTER_CMD_OPTION_LOCAL_ADDR_FIELD			(`NIF_MASTER_CMD_OPTION_LOCAL_ADDR_HIGH):(`NIF_MASTER_CMD_OPTION_LOCAL_ADDR_LOW)

// extended address 9-26-2014
`define NIF_MASTER_CMD_OPTION_EXT_ADDR_WIDTH			28
`define NIF_MASTER_CMD_OPTION_EXT_ADDR_LOW				(`NIF_MASTER_CMD_OPTION_LOCAL_ADDR_HIGH + 1)
`define NIF_MASTER_CMD_OPTION_EXT_ADDR_HIGH				(`NIF_MASTER_CMD_OPTION_EXT_ADDR_LOW + `NIF_MASTER_CMD_OPTION_EXT_ADDR_WIDTH - 1)
`define	NIF_MASTER_CMD_OPTION_EXT_ADDR_FIELD			(`NIF_MASTER_CMD_OPTION_EXT_ADDR_HIGH):(`NIF_MASTER_CMD_OPTION_EXT_ADDR_LOW)

`define NIF_MASTER_CMD_OPTION_ADDR_WIDTH				64
`define NIF_MASTER_CMD_OPTION_ADDR_LOW					(`NIF_MASTER_CMD_OPTION_LOCAL_ADDR_LOW)
`define NIF_MASTER_CMD_OPTION_ADDR_HIGH					(`NIF_MASTER_CMD_OPTION_ADDR_LOW + `NIF_MASTER_CMD_OPTION_ADDR_WIDTH - 1)
`define NIF_MASTER_CMD_OPTION_ADDR_FIELD				(`NIF_MASTER_CMD_OPTION_ADDR_HIGH):(`NIF_MASTER_CMD_OPTION_ADDR_LOW)

`define NIF_MASTER_CMD_OPTION_TRANSACTION_OPTIONS_WIDTH	4
`define	NIF_MASTER_CMD_OPTION_TRANSACTION_OPTIONS_LOW	(`NIF_MASTER_CMD_OPTION_EXT_ADDR_HIGH + 1)
`define NIF_MASTER_CMD_OPTION_TRANSACTION_OPTIONS_HIGH	(`NIF_MASTER_CMD_OPTION_TRANSACTION_OPTIONS_LOW + `NIF_MASTER_CMD_OPTION_TRANSACTION_OPTIONS_WIDTH - 1)
`define	NIF_MASTER_CMD_OPTION_TRANSACTION_OPTIONS_FIELD	(`NIF_MASTER_CMD_OPTION_TRANSACTION_OPTIONS_HIGH):(`NIF_MASTER_CMD_OPTION_TRANSACTION_OPTIONS_LOW)

`define	NIF_MASTER_CMD_OPTION_LOCAL_FLOW_WIDTH			10
`define	NIF_MASTER_CMD_OPTION_LOCAL_FLOW_LOW			(`NIF_MASTER_CMD_OPTION_TRANSACTION_OPTIONS_HIGH + 1)
`define	NIF_MASTER_CMD_OPTION_LOCAL_FLOW_HIGH			(`NIF_MASTER_CMD_OPTION_LOCAL_FLOW_LOW + `NIF_MASTER_CMD_OPTION_LOCAL_FLOW_WIDTH - 1)
`define	NIF_MASTER_CMD_OPTION_LOCAL_FLOW_FIELD			(`NIF_MASTER_CMD_OPTION_LOCAL_FLOW_HIGH):(`NIF_MASTER_CMD_OPTION_LOCAL_FLOW_LOW)



`define	NIF_MASTER_CMD_OPTION_RESERVED_WIDTH		10

//`define	NIF_MASTER_CMD_OPTION_WIDTH					(`NIF_MASTER_CMD_OPTION_LENGTH_WIDTH + `NIF_MASTER_CMD_OPTION_LOCAL_ADDR_WIDTH + `NIF_MASTER_CMD_OPTION_TRANSACTION_ID_WIDTH + `NIF_MASTER_CMD_OPTION_LOCAL_FLOW_WIDTH + `NIF_MASTER_CMD_OPTION_RESERVED_WIDTH + NIF_MASTER_CMD_OPTION_EXT_ADDR_WIDTH)

`define	NIF_MASTER_CMD_OPTION_WIDTH					(`NIF_MASTER_CMD_OPTION_LENGTH_WIDTH + `NIF_MASTER_CMD_OPTION_LOCAL_ADDR_WIDTH + `NIF_MASTER_CMD_OPTION_LOCAL_FLOW_WIDTH  + `NIF_MASTER_CMD_OPTION_EXT_ADDR_WIDTH + `NIF_MASTER_CMD_OPTION_TRANSACTION_OPTIONS_WIDTH)

////////////////////////////////////////
//}}} MASTER INTERFACE
////////////////////////////////////////



////////////////////////////////////////
//{{{ MESSAGE INTERFACE
////////////////////////////////////////

// ---------------------------------
// MSG HEADER FIELD DEFINITIONS
// ---------------------------------
`define	NIF_MSG_TYPE_WIDTH							8
`define	NIF_MSG_TYPE_LOW							0
`define	NIF_MSG_TYPE_HIGH							(`NIF_MSG_TYPE_LOW + `NIF_MSG_TYPE_WIDTH - 1)
`define	NIF_MSG_TYPE_FIELD							(`NIF_MSG_TYPE_HIGH):(`NIF_MSG_TYPE_LOW)
`define	NIF_MSG_TGT_DEVICE_ID_WIDTH					16
`define	NIF_MSG_TGT_DEVICE_ID_LOW					(`NIF_MSG_TYPE_HIGH + 1)
`define	NIF_MSG_TGT_DEVICE_ID_HIGH					(`NIF_MSG_TGT_DEVICE_ID_LOW + `NIF_MSG_TGT_DEVICE_ID_WIDTH - 1)
`define	NIF_MSG_TGT_DEVICE_ID_FIELD					(`NIF_MSG_TGT_DEVICE_ID_HIGH):(`NIF_MSG_TGT_DEVICE_ID_LOW)
`define	NIF_MSG_INIT_DEVICE_ID_WIDTH				16
`define	NIF_MSG_INIT_DEVICE_ID_LOW					(`NIF_MSG_TGT_DEVICE_ID_HIGH + 1)
`define	NIF_MSG_INIT_DEVICE_ID_HIGH					(`NIF_MSG_INIT_DEVICE_ID_LOW + `NIF_MSG_INIT_DEVICE_ID_WIDTH - 1)
`define	NIF_MSG_INIT_DEVICE_ID_FIELD				(`NIF_MSG_INIT_DEVICE_ID_HIGH):(`NIF_MSG_INIT_DEVICE_ID_LOW)
`define	NIF_MSG_LENGTH_WIDTH						10
`define	NIF_MSG_LENGTH_LOW							(`NIF_MSG_INIT_DEVICE_ID_HIGH + 1)
`define	NIF_MSG_LENGTH_HIGH							(`NIF_MSG_LENGTH_LOW + `NIF_MSG_LENGTH_WIDTH - 1)
`define	NIF_MSG_LENGTH_FIELD						(`NIF_MSG_LENGTH_HIGH):(`NIF_MSG_LENGTH_LOW)
`define	NIF_MSG_COMPLETION_REQUIRED_FLAG			(`NIF_MSG_LENGTH_HIGH + 1)
`define NIF_MSG_TRANSACTION_ID_WIDTH				10
`define NIF_MSG_TRANSACTION_ID_LOW					64
`define NIF_MSG_TRANSACTION_ID_HIGH					(`NIF_MSG_TRANSACTION_ID_LOW + `NIF_MSG_TRANSACTION_ID_WIDTH - 1)
`define NIF_MSG_TRANSACTION_ID_FIELD				(`NIF_MSG_TRANSACTION_ID_HIGH):(`NIF_MSG_TRANSACTION_ID_LOW)
`define NIF_MSG_ERROR_CODE_WIDTH					7
`define NIF_MSG_ERROR_CODE_LOW						80
`define NIF_MSG_ERROR_CODE_HIGH						(`NIF_MSG_ERROR_CODE_LOW + `NIF_MSG_ERROR_CODE_WIDTH - 1)
`define NIF_MSG_ERROR_CODE_FIELD					(`NIF_MSG_ERROR_CODE_HIGH):(`NIF_MSG_ERROR_CODE_LOW)
`define NIF_MSG_HEADER_RESERVED_WIDTH				(128-(`NIF_MSG_ERROR_CODE_HIGH + 1))
`define	NIF_MSG_HEADER_RESERVED_FIELD				(127):(`NIF_MSG_ERROR_CODE_HIGH + 1)
// MSG_LENGTH includes this 16 byte header
// Maximum message length including the header is 1008 bytes. (Maximum pure payload is 992 bytes)
// Message length must be multiple of 16 currently.


// ---------------------------------
// ERROR DEFINITIONS
// ---------------------------------
`define	NIF_MSG_SEND_ERROR_OKAY						2'd0
`define	NIF_MSG_SEND_ERROR_RETRY					2'd1
`define	NIF_MSG_SEND_ERROR_LOCAL_FATAL				2'd2
`define	NIF_MSG_SEND_ERROR_REMOTE_FATAL				2'd3


// ---------------------------------
// MESSAGE TYPE DEFINITIONS
// ---------------------------------
// 0x00 - 0x1F : Reserved for system messages
// 0x20 - 0x2F : Reserved for memory request commands
`define	NIF_MSG_TYPE_MEMORY_DMA_REQUEST				8'h20
`define	NIF_MSG_TYPE_MEMORY_DMA_COMPLETE			8'h21
`define SAP_MSG_TYPE_EXECUTE_REQUEST				8'h22
`define SAP_MSG_TYPE_EXECUTE_COMPLETE				8'h23
// 0x30 - 0xFF : Not yet reserved

////////////////////////////////////////
//}}} MESSAGE INTERFACE
////////////////////////////////////////



////////////////////////////////////////
//{{{ DMA DESCRIPTOR FIELD DEFINITIONS
////////////////////////////////////////

`define	NIF_DMA_DESCRIPTOR_LENGTH_WIDTH		36
`define	NIF_DMA_DESCRIPTOR_LENGTH_LOW		0
`define	NIF_DMA_DESCRIPTOR_LENGTH_HIGH		(`NIF_DMA_DESCRIPTOR_LENGTH_LOW + `NIF_DMA_DESCRIPTOR_LENGTH_WIDTH - 1)
`define	NIF_DMA_DESCRIPTOR_LENGTH_FIELD		(`NIF_DMA_DESCRIPTOR_LENGTH_HIGH):(`NIF_DMA_DESCRIPTOR_LENGTH_LOW)

`define	NIF_DMA_DESCRIPTOR_DEVICE_WIDTH		16
`define	NIF_DMA_DESCRIPTOR_DEVICE_LOW		(`NIF_DMA_DESCRIPTOR_LENGTH_HIGH + 1)
`define	NIF_DMA_DESCRIPTOR_DEVICE_HIGH		(`NIF_DMA_DESCRIPTOR_DEVICE_LOW + `NIF_DMA_DESCRIPTOR_DEVICE_WIDTH - 1)
`define	NIF_DMA_DESCRIPTOR_DEVICE_FIELD		(`NIF_DMA_DESCRIPTOR_DEVICE_HIGH):(`NIF_DMA_DESCRIPTOR_DEVICE_LOW)

`define	NIF_DMA_DESCRIPTOR_FLOW_WIDTH		10
`define	NIF_DMA_DESCRIPTOR_FLOW_LOW			(`NIF_DMA_DESCRIPTOR_DEVICE_HIGH + 1)
`define	NIF_DMA_DESCRIPTOR_FLOW_HIGH		(`NIF_DMA_DESCRIPTOR_FLOW_LOW + `NIF_DMA_DESCRIPTOR_FLOW_WIDTH - 1)
`define	NIF_DMA_DESCRIPTOR_FLOW_FIELD		(`NIF_DMA_DESCRIPTOR_FLOW_HIGH):(`NIF_DMA_DESCRIPTOR_FLOW_LOW)

`define	NIF_DMA_DESCRIPTOR_RSVD				(`NIF_DMA_DESCRIPTOR_FLOW_HIGH + 1)
`define	NIF_DMA_DESCRIPTOR_LAST_TARGET_FLAG	(`NIF_DMA_DESCRIPTOR_RSVD + 1)

`define	NIF_DMA_DESCRIPTOR_ADDRESS_WIDTH	64
`define	NIF_DMA_DESCRIPTOR_ADDRESS_LOW		(`NIF_DMA_DESCRIPTOR_LAST_TARGET_FLAG + 1)
`define	NIF_DMA_DESCRIPTOR_ADDRESS_HIGH		(`NIF_DMA_DESCRIPTOR_ADDRESS_LOW + `NIF_DMA_DESCRIPTOR_ADDRESS_WIDTH - 1)
`define	NIF_DMA_DESCRIPTOR_ADDRESS_FIELD	(`NIF_DMA_DESCRIPTOR_ADDRESS_HIGH):(`NIF_DMA_DESCRIPTOR_ADDRESS_LOW)

`define NIF_DMA_DESCRIPTOR_ADDRESS_EXT_WIDTH 64
////////////////////////////////////////
//}}} DMA DESCRIPTOR FIELD DEFINITIONS
////////////////////////////////////////



////////////////////////////////////////
//{{{ WINDOW DESCRIPTOR FIELD DEFINITIONS
////////////////////////////////////////

`define	NIF_WINDOW_DESCRIPTOR_BURST_SIZE_WIDTH		12
`define	NIF_WINDOW_DESCRIPTOR_BURST_SIZE_LOW		0
`define	NIF_WINDOW_DESCRIPTOR_BURST_SIZE_HIGH		(`NIF_WINDOW_DESCRIPTOR_BURST_SIZE_LOW + `NIF_WINDOW_DESCRIPTOR_BURST_SIZE_WIDTH - 1)
`define	NIF_WINDOW_DESCRIPTOR_BURST_SIZE_FIELD		(`NIF_WINDOW_DESCRIPTOR_BURST_SIZE_HIGH):(`NIF_WINDOW_DESCRIPTOR_BURST_SIZE_LOW)

`define	NIF_WINDOW_DESCRIPTOR_BURST_STRIDE_WIDTH	12
`define	NIF_WINDOW_DESCRIPTOR_BURST_STRIDE_LOW		(`NIF_WINDOW_DESCRIPTOR_BURST_SIZE_HIGH + 1)
`define	NIF_WINDOW_DESCRIPTOR_BURST_STRIDE_HIGH		(`NIF_WINDOW_DESCRIPTOR_BURST_STRIDE_LOW + `NIF_WINDOW_DESCRIPTOR_BURST_STRIDE_WIDTH - 1)
`define	NIF_WINDOW_DESCRIPTOR_BURST_STRIDE_FIELD	(`NIF_WINDOW_DESCRIPTOR_BURST_STRIDE_HIGH):(`NIF_WINDOW_DESCRIPTOR_BURST_STRIDE_LOW)

`define	NIF_WINDOW_DESCRIPTOR_NUM_BURST_WIDTH		11
`define	NIF_WINDOW_DESCRIPTOR_NUM_BURST_LOW			(`NIF_WINDOW_DESCRIPTOR_BURST_STRIDE_HIGH + 1)
`define	NIF_WINDOW_DESCRIPTOR_NUM_BURST_HIGH		(`NIF_WINDOW_DESCRIPTOR_NUM_BURST_LOW + `NIF_WINDOW_DESCRIPTOR_NUM_BURST_WIDTH - 1)
`define	NIF_WINDOW_DESCRIPTOR_NUM_BURST_FIELD		(`NIF_WINDOW_DESCRIPTOR_NUM_BURST_HIGH):(`NIF_WINDOW_DESCRIPTOR_NUM_BURST_LOW)

`define	NIF_WINDOW_DESCRIPTOR_VALID_FLAG			(`NIF_WINDOW_DESCRIPTOR_NUM_BURST_HIGH + 1)

////////////////////////////////////////
//}}} WINDOW DESCRIPTOR FIELD DEFINITIONS
////////////////////////////////////////
