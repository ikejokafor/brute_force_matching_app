`include "math.vh"

`define AXH_CTAG_WIDTH 						8
`define AXH_CTAGPAR_WIDTH 					1
`define AXH_COM_WIDTH 						13
`define AXH_COMPAR_WIDTH					1
`define AXH_CABT_WIDTH						3
`define AXH_CEA_WIDTH						64
`define AXH_CEAPAR_WIDTH					1
`define AXH_CCH_WIDTH						16
`define AXH_CSIZE_WIDTH						12
`define AXH_CROOM_WIDTH						8

`define MAX_NUM_OUTSTANDING_COMMANDS 		32
`define MAX_NUM_TAGS 						`MAX_NUM_OUTSTANDING_COMMANDS
`define TAG_WIDTH 							clog2(`MAX_NUM_OUTSTANDING_COMMANDS)

`define	INTERRUPT_SOURCE_WIDTH				11

`define READ_CL_S							13'h0A50
`define READ_CL_M							13'h0A60
`define READ_CL_LCK							13'h0A6B
`define READ_CL_RES							13'h0A67
`define TOUCH_I								13'h0240
`define TOUCH_S								13'h0250
`define TOUCH_M								13'h0260
`define WRITE_MI							13'h0D60
`define WRITE_MS							13'h0D70
`define WRITE_UNLOCK						13'h0D6B
`define WRITE_C								13'h0D67
`define PUSH_I								13'h0140
`define PUSH_S								13'h0150
`define EVICT_I								13'h1140
`define ZERO_M								13'h1260
`define LOCK								13'h016B
`define UNLOCK								13'h017B
`define READ_CL_NA							13'h0A00
`define READ_PNA							13'h0E00
`define WRITE_NA							13'h0D00
`define WRITE_INJ							13'h0D10
`define FLUSH								13'h0100
`define INTREQ								13'h0000
`define RESTART								13'h0001
`define RESTART_ODD_PARITY					1
`define RESTART_EVEN_PARITY					0

`define COMMAND_ARRAY_CTAG_LOW				0
`define COMMAND_ARRAY_CTAG_HIGH				(`COMMAND_ARRAY_CTAG_LOW + `AXH_CTAG_WIDTH - 1)
`define COMMAND_ARRAY_CTAG_FIELD			(`COMMAND_ARRAY_CTAG_HIGH):(`COMMAND_ARRAY_CTAG_LOW)
`define COMMAND_ARRAY_CEA_LOW				(`COMMAND_ARRAY_CTAG_HIGH + 1)
`define COMMAND_ARRAY_CEA_HIGH				(`COMMAND_ARRAY_CEA_LOW + `AXH_CEA_WIDTH - 1)
`define COMMAND_ARRAY_CEA_FIELD				(`COMMAND_ARRAY_CEA_HIGH):(`COMMAND_ARRAY_CEA_LOW)
`define COMMAND_ARRAY_COM_LOW				(`COMMAND_ARRAY_CEA_HIGH + 1)
`define COMMAND_ARRAY_COM_HIGH				(`COMMAND_ARRAY_COM_LOW + `AXH_COM_WIDTH - 1)
`define COMMAND_ARRAY_COM_FIELD				(`COMMAND_ARRAY_COM_HIGH):(`COMMAND_ARRAY_COM_LOW)
`define COMMAND_ARRAY_CSIZE_LOW				(`COMMAND_ARRAY_COM_HIGH + 1)
`define COMMAND_ARRAY_CSIZE_HIGH			(`COMMAND_ARRAY_CSIZE_LOW + `AXH_CSIZE_WIDTH - 1)
`define COMMAND_ARRAY_CSIZE_FIELD			(`COMMAND_ARRAY_CSIZE_HIGH):(`COMMAND_ARRAY_CSIZE_LOW)
`define COMMAND_ARRAY_CABT_LOW				(`COMMAND_ARRAY_CSIZE_HIGH + 1)
`define COMMAND_ARRAY_CABT_HIGH				(`COMMAND_ARRAY_CABT_LOW + `AXH_CABT_WIDTH - 1)
`define COMMAND_ARRAY_CABT_FIELD			(`COMMAND_ARRAY_CABT_HIGH):(`COMMAND_ARRAY_CABT_LOW)
`define COMMAND_ARRAY_CCH_LOW				(`COMMAND_ARRAY_CABT_HIGH + 1)
`define COMMAND_ARRAY_CCH_HIGH				(`COMMAND_ARRAY_CCH_LOW + `AXH_CCH_WIDTH - 1)
`define COMMAND_ARRAY_CCH_FIELD				(`COMMAND_ARRAY_CCH_HIGH):(`COMMAND_ARRAY_CCH_LOW)
`define COMMAND_ARRAY_CTAGPAR_FLAG			(`COMMAND_ARRAY_CCH_HIGH + 1)
`define COMMAND_ARRAY_CEAPAR_FLAG			(`COMMAND_ARRAY_CTAGPAR_FLAG + 1)
`define COMMAND_ARRAY_COMPAR_FLAG			(`COMMAND_ARRAY_CEAPAR_FLAG + 1)

`define COMMAND_ORDERING_STRICT				3'b000
`define COMMAND_ORDERING_ABORT				3'b001
`define COMMAND_ORDERING_PAGE				3'b010
`define COMMAND_ORDERING_PREF				3'b011
`define COMMAND_ORDERING_SPEC				3'b111

`define	COMMAND_STATE_IDLE		    		3'b000
`define	COMMAND_STATE_PENDING      			3'b001
`define	COMMAND_STATE_ISSUED      			3'b010
`define	COMMAND_STATE_FLUSHED      			3'b011
`define	COMMAND_STATE_RESTART_REQUEST		3'b100
`define	COMMAND_STATE_RESTART_PENDING		3'b101
`define	COMMAND_STATE_RESTART_REISSUE		3'b110
`define	COMMAND_STATE_COMPLETE      		3'b111
`define COMMAND_STATE_WIDTH 				3

`define RESPONSE_DONE						8'h00
`define RESPONSE_AERROR						8'h01
`define RESPONSE_DERROR						8'h03
`define RESPONSE_NLOCK						8'h04
`define RESPONSE_NRES						8'h05
`define RESPONSE_FLUSHED					8'h06
`define RESPONSE_FAULT						8'h07
`define RESPONSE_FAILED						8'h08
`define RESPONSE_PAGED						8'h0A

`define PSL_CONTROL_START					8'h90
`define PSL_CONTROL_RESET					8'h80
`define PSL_CONTROL_TIMEBASE				8'h42

`define TRANSACTION_INFO_COMMAND_WIDTH		`AXH_COM_WIDTH
`define TRANSACTION_INFO_COMMAND_LOW		0
`define TRANSACTION_INFO_COMMAND_HIGH		(`TRANSACTION_INFO_COMMAND_LOW + `TRANSACTION_INFO_COMMAND_WIDTH - 1)
`define TRANSACTION_INFO_COMMAND_FIELD  	(`TRANSACTION_INFO_COMMAND_HIGH):(`TRANSACTION_INFO_COMMAND_LOW)
`define TRANSACTION_INFO_TAG_WIDTH			`TAG_WIDTH
`define TRANSACTION_INFO_TAG_LOW			(`TRANSACTION_INFO_COMMAND_HIGH + 1)
`define TRANSACTION_INFO_TAG_HIGH			(`TRANSACTION_INFO_TAG_LOW + `TRANSACTION_INFO_TAG_WIDTH - 1)
`define TRANSACTION_INFO_TAG_FIELD			(`TRANSACTION_INFO_TAG_HIGH):(`TRANSACTION_INFO_TAG_LOW)
`define TRANSACTION_INFO_LENGTH_WIDTH		13
`define TRANSACTION_INFO_LENGTH_LOW			(`TRANSACTION_INFO_TAG_HIGH + 1)
`define TRANSACTION_INFO_LENGTH_HIGH		(`TRANSACTION_INFO_LENGTH_LOW + `TRANSACTION_INFO_LENGTH_WIDTH - 1)
`define TRANSACTION_INFO_LENGTH_FIELD		(`TRANSACTION_INFO_LENGTH_HIGH):(`TRANSACTION_INFO_LENGTH_LOW)
`define TRANSACTION_INFO_OFFSET_WIDTH		8
`define TRANSACTION_INFO_OFFSET_LOW			(`TRANSACTION_INFO_LENGTH_HIGH + 1)
`define TRANSACTION_INFO_OFFSET_HIGH		(`TRANSACTION_INFO_OFFSET_LOW + `TRANSACTION_INFO_OFFSET_WIDTH - 1)
`define TRANSACTION_INFO_OFFSET_FIELD		(`TRANSACTION_INFO_OFFSET_HIGH):(`TRANSACTION_INFO_OFFSET_LOW)
`define TRANSACTION_INFO_ADDRESS_WIDTH		64
`define TRANSACTION_INFO_ADDRESS_LOW		(`TRANSACTION_INFO_OFFSET_HIGH + 1)
`define TRANSACTION_INFO_ADDRESS_HIGH		(`TRANSACTION_INFO_ADDRESS_LOW + `TRANSACTION_INFO_ADDRESS_WIDTH - 1)
`define TRANSACTION_INFO_ADDRESS_FIELD		(`TRANSACTION_INFO_ADDRESS_HIGH):(`TRANSACTION_INFO_ADDRESS_LOW)
`define TRANSACTION_INFO_SOURCE_WIDTH		3
`define TRANSACTION_INFO_SOURCE_LOW			(`TRANSACTION_INFO_ADDRESS_HIGH + 1)
`define TRANSACTION_INFO_SOURCE_HIGH		(`TRANSACTION_INFO_SOURCE_LOW + `TRANSACTION_INFO_SOURCE_WIDTH - 1)
`define TRANSACTION_INFO_SOURCE_FIELD		(`TRANSACTION_INFO_SOURCE_HIGH):(`TRANSACTION_INFO_SOURCE_LOW)
`define TRANSACTION_INFO_RNW_WIDTH			1
`define TRANSACTION_INFO_RNW_LOW			(`TRANSACTION_INFO_SOURCE_HIGH + 1)
`define TRANSACTION_INFO_RNW_HIGH			(`TRANSACTION_INFO_RNW_LOW + `TRANSACTION_INFO_RNW_WIDTH - 1)
`define TRANSACTION_INFO_RNW_FIELD			(`TRANSACTION_INFO_RNW_HIGH):(`TRANSACTION_INFO_RNW_LOW)
`define TRANSACTION_INFO_WIDTH				(`TRANSACTION_INFO_COMMAND_WIDTH + `TRANSACTION_INFO_TAG_WIDTH + `TRANSACTION_INFO_LENGTH_WIDTH + `TRANSACTION_INFO_OFFSET_WIDTH + `TRANSACTION_INFO_ADDRESS_WIDTH + `TRANSACTION_INFO_SOURCE_WIDTH + `TRANSACTION_INFO_RNW_WIDTH)
`define TRANSACTION_INFO_LOW				0
`define TRANSACTION_INFO_HIGH				(`TRANSACTION_INFO_LOW + `TRANSACTION_INFO_WIDTH - 1)
`define TRANSACTION_INFO_FIELD				(`TRANSACTION_INFO_HIGH):(`TRANSACTION_INFO_LOW)

`define READ_INFO_OFFSET_WIDTH				8
`define READ_INFO_OFFSET_LOW				0
`define READ_INFO_OFFSET_HIGH				(`READ_INFO_OFFSET_LOW + `READ_INFO_OFFSET_WIDTH - 1)
`define READ_INFO_OFFSET_FIELD				(`READ_INFO_OFFSET_HIGH):(`READ_INFO_OFFSET_LOW)
`define READ_INFO_LENGTH_WIDTH				8
`define READ_INFO_LENGTH_LOW				(`READ_INFO_OFFSET_HIGH + 1)
`define READ_INFO_LENGTH_HIGH				(`READ_INFO_LENGTH_LOW + `READ_INFO_LENGTH_WIDTH - 1)
`define READ_INFO_LENGTH_FIELD				(`READ_INFO_LENGTH_HIGH):(`READ_INFO_LENGTH_LOW)
`define READ_INFO_TAG_WIDTH					5
`define READ_INFO_TAG_LOW					(`READ_INFO_LENGTH_HIGH + 1)
`define READ_INFO_TAG_HIGH					(`READ_INFO_TAG_LOW + `READ_INFO_TAG_WIDTH - 1)
`define READ_INFO_TAG_FIELD					(`READ_INFO_TAG_HIGH):(`READ_INFO_TAG_LOW)

`define WRITE_INFO_OFFSET_WIDTH				8
`define WRITE_INFO_OFFSET_LOW				0
`define WRITE_INFO_OFFSET_HIGH				(`WRITE_INFO_OFFSET_LOW + `WRITE_INFO_OFFSET_WIDTH - 1)
`define WRITE_INFO_OFFSET_FIELD				(`WRITE_INFO_OFFSET_HIGH):(`WRITE_INFO_OFFSET_LOW)
`define WRITE_INFO_LENGTH_WIDTH				8
`define WRITE_INFO_LENGTH_LOW				(`WRITE_INFO_OFFSET_HIGH + 1)
`define WRITE_INFO_LENGTH_HIGH				(`WRITE_INFO_LENGTH_LOW + `WRITE_INFO_LENGTH_WIDTH - 1)
`define WRITE_INFO_LENGTH_FIELD				(`WRITE_INFO_LENGTH_HIGH):(`WRITE_INFO_LENGTH_LOW)
`define WRITE_INFO_TAG_WIDTH				5
`define WRITE_INFO_TAG_LOW					(`WRITE_INFO_LENGTH_HIGH + 1)
`define WRITE_INFO_TAG_HIGH					(`WRITE_INFO_TAG_LOW + `WRITE_INFO_TAG_WIDTH - 1)
`define WRITE_INFO_TAG_FIELD				(`WRITE_INFO_TAG_HIGH):(`WRITE_INFO_TAG_LOW)
`define WRITE_INFO_BUFFER_ADV_FLAG_WIDTH	1
`define WRITE_INFO_BUFFER_ADV_FLAG_LOW		(`WRITE_INFO_TAG_HIGH + 1)
`define WRITE_INFO_BUFFER_ADV_FLAG_HIGH		(`WRITE_INFO_BUFFER_ADV_FLAG_LOW + `WRITE_INFO_BUFFER_ADV_FLAG_WIDTH - 1)
`define WRITE_INFO_BUFFER_ADV_FLAG			(`WRITE_INFO_BUFFER_ADV_FLAG_HIGH):(`WRITE_INFO_BUFFER_ADV_FLAG_LOW)

`define INTERRUPT_INFO_SOURCE_WIDTH			`INTERRUPT_SOURCE_WIDTH
`define INTERRUPT_INFO_SOURCE_LOW			0
`define INTERRUPT_INFO_SOURCE_HIGH			(`INTERRUPT_INFO_SOURCE_LOW + `INTERRUPT_INFO_SOURCE_WIDTH - 1)
`define INTERRUPT_INFO_SOURCE_FIELD			(`INTERRUPT_INFO_SOURCE_HIGH):(`INTERRUPT_INFO_SOURCE_LOW)
`define INTERRUPT_INFO_TAG_WIDTH			5
`define INTERRUPT_INFO_TAG_LOW				(`INTERRUPT_INFO_SOURCE_HIGH + 1)
`define INTERRUPT_INFO_TAG_HIGH				(`INTERRUPT_INFO_TAG_LOW + `INTERRUPT_INFO_TAG_WIDTH - 1)
`define INTERRUPT_INFO_TAG_FIELD			(`INTERRUPT_INFO_TAG_HIGH):(`INTERRUPT_INFO_TAG_LOW)

`define READ_INFO_WIDTH 					(`READ_INFO_OFFSET_WIDTH + `READ_INFO_LENGTH_WIDTH + `READ_INFO_TAG_WIDTH)
`define WRITE_INFO_WIDTH 					(`WRITE_INFO_OFFSET_WIDTH + `WRITE_INFO_LENGTH_WIDTH + `WRITE_INFO_TAG_WIDTH + `WRITE_INFO_BUFFER_ADV_FLAG_WIDTH)
`define INTERRUPT_INFO_WIDTH				(`INTERRUPT_INFO_SOURCE_WIDTH + `INTERRUPT_INFO_TAG_WIDTH)

`define STATE_VECTOR_WIDTH					(`MAX_NUM_OUTSTANDING_COMMANDS*`COMMAND_STATE_WIDTH)
`define COMMAND_WIDTH 						(`AXH_CSIZE_WIDTH + `AXH_COM_WIDTH + `AXH_CTAG_WIDTH + `AXH_CEA_WIDTH + `AXH_CABT_WIDTH + `AXH_CCH_WIDTH + `AXH_CTAGPAR_WIDTH + `AXH_CEAPAR_WIDTH + `AXH_COMPAR_WIDTH)
`define CACHELINE_SIZE_BYTES				128

